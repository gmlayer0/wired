// top level of dcache