// 此文件是核心的顶层
`include "wired0_defines.svh"

module wired_top(
    `_WIRED_GENERAL_DEFINE
);

endmodule