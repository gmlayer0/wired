// Wired2 下一代缓存模块
// 这个模块只负责进行缓存命中判断，永不阻塞
