`include "tl_util.svh"

module wired_mp #(
  parameter int CPU_NUM = 4
) (
  input clk,
  input rst_n
);

endmodule
