`ifndef _WIRED_HEADER
`define _WIRED_HEADER

`define _VERILATOR
// `define _ASIC

`include "wired0_params.svh"
`include "wired0_decoder.svh"
`include "wired0_macros.svh"
`include "wired0_structure.svh"
`include "wired0_csr.svh"

`endif
