`ifndef _WIRED_HEADER
`define _WIRED_HEADER

`include "wired0_structure.svh"
`include "wired0_macros.svh"

`endif
