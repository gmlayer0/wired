// Wired2 乱序访存模块 wired_lsung
// ng means Next Gen

// 该模块内建一个非阻塞缓存，

`include "wired0_defines.svh"

module wired_lsung(

);

endmodule
