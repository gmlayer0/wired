`ifndef _WIRED_HEADER
`define _WIRED_HEADER

`include "wired0_decoder.svh"
`include "wired0_macros.svh"
`include "wired0_params.svh"
`include "wired0_structure.svh"

`endif
